module IFU (
	input clk,
	input rst,
	input [`XLEN-1:0] pc,
	output [31:0] inst
);

	//assign inst = pmem_read[pc];

endmodule //IFU