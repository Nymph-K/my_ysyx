module ex_mem_reg (
    input           clk                 ,
    input           rst                 ,

    input           mem_idle            ,
    input           in_valid            ,
    input           in_ready            ,
    input  [ 2:0]   in_funct3           ,
    input  [31:0]   in_pc               ,
    input  [31:0]   in_inst             ,
    input  [ 4:0]   in_rs1              ,
    input  [ 4:0]   in_rs2              ,
    input  [63:0]   in_x_rs2            ,
    input  [63:0]   in_x_rd             ,
    input  [ 4:0]   in_rd               ,
    input           in_rd_idx_0         ,
    input           in_rd_w_en          ,
    input           in_rd_w_src_exu     ,
    input           in_rd_w_src_mem     ,
    input           in_rd_w_src_csr     ,
    input           in_csr_w_en         ,
    input  [11:0]   in_csr_addr         ,
    input  [63:0]   in_csr_r_data       ,
    input  [63:0]   in_exu_result       ,
    input           in_inst_system_ebreak,
    input           in_inst_load        ,
    input           in_inst_store       ,

    output reg          out_valid           ,
    output              out_ready           ,
    output reg [ 2:0]   out_funct3          ,
    output reg [31:0]   out_pc              ,
    output reg [31:0]   out_inst            ,
    output reg [ 4:0]   out_rs1             ,
    output reg [ 4:0]   out_rs2             ,
    output reg [63:0]   out_x_rs2           ,
    output reg [63:0]   out_x_rd            ,
    output reg [ 4:0]   out_rd              ,
    output reg          out_rd_idx_0        ,
    output reg          out_rd_w_en         ,
    output reg          out_rd_w_src_exu    ,
    output reg          out_rd_w_src_mem    ,
    output reg          out_rd_w_src_csr    ,
    output reg          out_csr_w_en        ,
    output reg [11:0]   out_csr_addr        ,
    output reg [63:0]   out_csr_r_data      ,
    output reg [63:0]   out_exu_result      ,
    output reg          out_inst_system_ebreak,
    output reg          out_inst_load       ,
    output reg          out_inst_store      
);

    wire stall = (~in_ready & out_valid) | ~mem_idle;
    wire wen = in_valid & ~stall;
    wire ctrl_flush = rst | (~in_valid & ~stall);
    assign out_ready = mem_idle & !(in_valid & ~in_ready & out_valid);
    
    always @(posedge clk ) begin
        if (ctrl_flush) begin
            out_valid               <= 0;
            out_rd_w_en             <= 0;
            out_csr_w_en            <= 0;
            out_inst_system_ebreak  <= 0;
            out_inst_load           <= 0;
            out_inst_store          <= 0;
        end else begin
            if(wen) begin
                out_valid               <= in_valid;
                out_rd_w_en             <= in_rd_w_en;
                out_csr_w_en            <= in_csr_w_en;
                out_inst_system_ebreak  <= in_inst_system_ebreak;
                out_inst_load           <= in_inst_load;
                out_inst_store          <= in_inst_store;
            end
        end
    end
    
    always @(posedge clk ) begin
        if (rst) begin
            out_funct3          <= 0;
            out_pc              <= 0;
            out_inst            <= 0;
            out_rs1             <= 0;
            out_rs2             <= 0;
            out_x_rs2           <= 0;
            out_x_rd            <= 0;
            out_rd              <= 0;
            out_rd_idx_0        <= 0;
            out_rd_w_src_exu    <= 0;
            out_rd_w_src_mem    <= 0;
            out_rd_w_src_csr    <= 0;
            out_csr_addr        <= 0;
            out_csr_r_data      <= 0;
            out_exu_result      <= 0;
        end else begin
            if(wen) begin
                out_funct3          <= in_funct3; 
                out_pc              <= in_pc; 
                out_inst            <= in_inst; 
                out_rs1             <= in_rs1; 
                out_rs2             <= in_rs2; 
                out_x_rs2           <= in_x_rs2; 
                out_x_rd            <= in_x_rd; 
                out_rd              <= in_rd; 
                out_rd_idx_0        <= in_rd_idx_0; 
                out_rd_w_src_exu    <= in_rd_w_src_exu; 
                out_rd_w_src_mem    <= in_rd_w_src_mem; 
                out_rd_w_src_csr    <= in_rd_w_src_csr; 
                out_csr_addr        <= in_csr_addr; 
                out_csr_r_data      <= in_csr_r_data; 
                out_exu_result      <= in_exu_result; 
            end
        end
    end

endmodule //ex_mem_reg
